library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity midori_roundconstants_enc is
	Port(
		i : in STD_LOGIC_VECTOR(4 downto 0); 
		o : out STD_LOGIC_VECTOR(127 downto 0)
	);
end midori_roundconstants_enc ;

architecture behavior of midori_roundconstants_enc is

type table is array (0 to 19) of STD_LOGIC_VECTOR(127 downto 0);

constant round_constants_enc : table := (
X"00000001000100010100010100000101",
X"00010101010000000101000000000000",
X"01000100000100000000010100010001",
X"00010100000001000000000100000101",
X"00000001000000000001000001010101",
X"01010001000000010001010100000000",
X"00000000000001000001010000010100",
X"00000000010001010101000001010000",
X"01000001000100000100000000000001",
X"00010000000000000100010101000000",
X"00010101000000010100000100010101",
X"00000100000001000100000001010100",
X"00010001000000010000010100000000",
X"01010101010000000101000001000100",
X"01010001010101010100000100000000",
X"00010101010100000100000000000001",
X"00000001010100000000010000010000",
X"00000100000001010100010100010000",
X"00010100000001000100000001000100",
X"00000000000000000000000000000000"
);

begin 

o <= round_constants_enc(to_integer(unsigned(i)));

end;

